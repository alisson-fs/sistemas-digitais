PACKAGE constants IS
  CONSTANT n : INTEGER := 4;
END PACKAGE constants;

