PACKAGE constants IS
	CONSTANT size : INTEGER := 4;
END PACKAGE constants;