PACKAGE constants IS
  CONSTANT n : INTEGER := 8;
END PACKAGE constants;